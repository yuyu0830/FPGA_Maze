library verilog;
use verilog.vl_types.all;
entity Top_tb is
end Top_tb;
