// parameter
parameter
    IDLE        = 3'b000,
    RUNNING     = 3'b001,
    MOVE        = 3'b010,
    LV_CHECK    = 3'b011,
    CLEAR       = 3'b100;

parameter
    PIXEL_EZ = 6'd40,
    PIXEL_MI = 6'd20,
    PIXEL_HD = 6'd16;

parameter
    ROW     = 6'd40,
    COLUMN  = 5'd30;

parameter
    LEFT    = 2'b00,
    UP      = 2'b01,
    DOWN    = 2'b10,
    RIGHT   = 2'b11;

parameter
    BLOCK_EZ_COL = 6'd16, // Eazy
    BLOCK_EZ_ROW = 5'd12,
    BLOCK_MI_COL = 6'd32, // Middle 
    BLOCK_MI_ROW = 5'd24,
    BLOCK_HD_COL = 6'd40, // Hard
    BLOCK_HD_ROW = 5'd30;

parameter
    [ROW * COLUMN - 1:0] MAZE_EZ = {
        40'b1111111111111111000000000000000000000000,
        40'b1010000000000001000000000000000000000000,
        40'b1010101111111101000000000000000000000000,
        40'b1000100010000001000000000000000000000000,
        40'b1110111010010111000000000000000000000000, // 5
        40'b1000100011110001000000000000000000000000,
        40'b1011101110000101000000000000000000000000,
        40'b1000001011110111000000000000000000000000,
        40'b1011101000000001000000000000000000000000,
        40'b1010101111011101000000000000000000000000, // 10
        40'b1000100001000101000000000000000000000000,
        40'b1111111111111111000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000, // 15
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000, // 20
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000, // 25
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000 // 30
    },
    MAZE_MI = {
        40'b1111111111111111111111111111111100000000,
        40'b1000001000000000000100000000000100000000,
        40'b1011101011111111110111011111110100000000,
        40'b1010001000001000010000010001000100000000,
        40'b1011101110101101011111111101011100000000, // 5
        40'b1000100010100101000000000001000100000000,
        40'b1010111011110101111111011111110100000000,
        40'b1010001000000101010000010000010100000000,
        40'b1011101110101101010111110111010100000000,
        40'b1000101010100101000001000100000100000000, // 10
        40'b1111101010101001110111011101111100000000,
        40'b1000001000101010010100000101000100000000,
        40'b1011111110111011010101110101110100000000,
        40'b1000000010000010010101000101000100000000,
        40'b1011111011111110110101011101011100000000, // 15
        40'b1000001000000010100101000100010100000000,
        40'b1011101110111010111101111111010100000000,
        40'b1010000010001000100101000001000100000000,
        40'b1010111111101110101101011101110100000000,
        40'b1010101000111010101111010101011100000000, // 20
        40'b1010001010000010101000010001000100000000,
        40'b1011101010111011101011011011010100000000,
        40'b1000100010001000000001001000010100000000,
        40'b1111111111111111111111111111111100000000,
        40'b0000000000000000000000000000000000000000, // 25
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000,
        40'b0000000000000000000000000000000000000000 // 30
    },
    MAZE_HD = {
        40'b1111111111111111111111111111111111111111,
        40'b1000001000000000010000000001000100000001,
        40'b1110101011101111011011110101011101010101,
        40'b1000100010001010001000010100000101010101,
        40'b1011111111101000100011011111111101011101,
        40'b1000000001000101010101000000000001010001,
        40'b1111111101111101011101111111111111010111,
        40'b1000000000000101000001000000010001010001,
        40'b1011111111111101011111110101110101011111,
        40'b1000100000010001010000010100000100000001,
        40'b1110101111010111110111010111111111111111,
        40'b1000100000100100010001000000000000000001,
        40'b1011101010111101011101111111111111111101,
        40'b1010001010000001000101010000000100000001,
        40'b1011111011111111110111010111110101111111,
        40'b1010000010000001000001000100010100000001,
        40'b1010111110111101011101011101110111111101,
        40'b1010101000100101010001110001010000000101,
        40'b1000001010001001011100000101000101110001,
        40'b1011111011111011010101111101111101010111,
        40'b1010000010000000000101000000000000010001,
        40'b1010111110111111111101111111111111111101,
        40'b1000100010100000000100010000000000000101,
        40'b1111101110111101111111010111111111011101,
        40'b1000100010000100000001000100000001000001,
        40'b1010101011110111110101111111011101111111,
        40'b1010001000010000000100010001010001000001,
        40'b1011111110111111111111010101110111011101,
        40'b1000000010000000000000000100000000000101,
        40'b1111111111111111111111111111111111111111
    };

