// parameter
parameter
    IDLE        = 3'b000,
    RUNNING     = 3'b001,
    MOVE        = 3'b010,
    LV_CHECK    = 3'b011,
    CLEAR       = 3'b100;

parameter
    ROW     = 7'd40,
    COLUMN  = 6'd30;

parameter
    LEFT    = 2'b00,
    UP      = 2'b01,
    DOWN    = 2'b10,
    RIGHT   = 2'b11;

parameter
    BLOCK_EZ_COL = 7'b16, // Eazy
    BLOCK_EZ_ROW = 6'b12,
    BLOCK_MI_COL = 7'b32, // Middle 
    BLOCK_MI_ROW = 6'b24,
    BLOCK_HD_COL = 7'b40, // Hard
    BLOCK_HD_ROW = 6'b30;

parameter
    [ROW * COLUMN:0] MAZE_EZ = {
        40'b10111_11111_11111_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000, // 5
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000, // 10
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b10000_00000_00000_10000_00000_00000_00000_00000,
        40'b11111_11111_11111_10000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000, // 15
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000, // 20
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000, // 25
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000 // 30
    },
    [ROW * COLUMN:0] MAZE_MI = {
        40'b10111_11111_11111_11111_11111_11000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000, // 5
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000, // 10
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000, // 15
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000, // 20
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b10000_00000_00000_00000_00000_01000_00000_00000,
        40'b11111_11111_11111_11111_11111_11000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000, // 25
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000,
        40'b00000_00000_00000_00000_00000_00000_00000_00000 // 30
    },
    [ROW * COLUMN:0] MAZE_HD = {
        40'b10111_11111_11111_11111_11111_11111_11111_11111,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001, // 5
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001, // 10
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001, // 15
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001, // 20
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001, // 25
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b10000_00000_00000_00000_00000_00000_00000_00001,
        40'b11111_11111_11111_11111_11111_11111_11111_11111 // 30
    };